package pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "./transaction_in.sv"
  `include "./transaction_out.sv"
  `include "./sequence_in.sv"

  `include "./sequencer.sv"
  `include "./driver.sv"
  `include "./monitor.sv"
  `include "./agent.sv"

  `include "./coverage.sv"
  `include "./scoreboard.sv"
  `include "./env.sv"
  `include "./simple_test.sv"
endpackage
